module mux_2to1(input [1:0]in,input select,output out);

    wire a1,a2;
    wire n_s;

    
    
endmodule