`include "mux_2to1.v"
module mux_4to1(input [3:0] in,input [1:0] select,output out);
    wire [1:0] m;

    
endmodule